Guitar mid scoop circuit

VIN 1 0 AC 300m
RIN 1 2 4.5k

RTPOT 2 20 150k
CTPOT 20 0 22u

RVOL1 2 3 0
RVOL2 3 0 250k

RMS 2 40 2.2k
*LMS 40 50 300m
LMS1 40 41 100m
LMS2 41 42 100m
LMS3 42 50 100m
K1 LMS1 LMS2 0.1
K2 LMS2 LMS3 0.1
K3 LMS1 LMS3 0.03
CMS 50 0 10n

.AC DEC 100 80 22000
.PLOT AC VDB(3) VP(3)

.END
